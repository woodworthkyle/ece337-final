library verilog;
use verilog.vl_types.all;
entity tb_memcontrol is
end tb_memcontrol;

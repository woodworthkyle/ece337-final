// $Id: $
// File name:   tb_mt48lc4m32b2
// Created:     12/4/2014
// Author:      Kyle Woodworth
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Testbench for SDRAM module

module tb_mt48lc4m32b2();
  
  initial begin
    
  end
  
endmodule
